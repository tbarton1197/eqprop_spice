.title testNetlist 
.SUBCKT neuron in out 
E1 2 0 in 0 4 
V1 out 2 0
F1 in 0 V1 0.25
X1 in 0 1N4148
X2 0 in 1N4148

.ENDS
.SUBCKT 1N4148 1 2 

R1 1 2 5.827E+9 
D1 1 2 1N4148
*
.MODEL 1N4148 D 
+ IS = 4.352E-9 
+ N = 1.906 
+ BV = 110 
+ IBV = 0.0001 
+ RS = 0.6458 
+ CJO = 7.048E-13 
+ VJ = 0.869 
+ M = 0.03 
+ FC = 0.5 
+ TT = 3.48E-9 
.ENDS
r_X1_in_00 X1_Nin_0 X1_in_0 420.0
r_X1_in_01 X1_Nin_1 X1_in_0 10.0
r_X1_in_10 X1_Nin_0 X1_in_1 420.0
r_X1_in_11 X1_Nin_1 X1_in_1 10.0
X1_neuron_0 X1_Nin_0 X2_in_0 neuron
X1_neuron_1 X1_Nin_1 X2_in_1 neuron
r_X2_in_00 output_net_0 X2_in_0 730.0
r_X2_in_01 output_net_1 X2_in_0 310.0
r_X2_in_10 output_net_0 X2_in_1 730.0
r_X2_in_11 output_net_1 X2_in_1 310.0
vin_0 X1_in_0 0 1
vin_1 X1_in_1 0 0
.op
.end
